/*---------------------------------------------------------------------------------------------------------
Name		:tb_tmds_encoder.v
Author		:Sesha Sayana Reddy Koppula
Student ID	:018399576
Description	:Test Bench for tmds_encoder.v
----------------------------------------------------------------------------------------------------------*/

`timescale 1ns/1ps

module tb_tmds_encoder;

    localparam integer C_PIXEL_DATA_WIDTH = 8;

    // Clocks & reset
    reg tmds_clk;   // 10x pixel clock
    reg pixel_clk;  // 1x pixel clock
    reg rst_n;

    // Pixel data
    reg [C_PIXEL_DATA_WIDTH-1:0] in_data_ch0; // Blue
    reg [C_PIXEL_DATA_WIDTH-1:0] in_data_ch1; // Green
    reg [C_PIXEL_DATA_WIDTH-1:0] in_data_ch2; // Red

    // Sync & DE
    reg hsync_pix_clk;
    reg vsync_pix_clk;
    reg de_pix_clk;

    // Outputs
    wire tmds_ch0_p, tmds_ch0_n;
    wire tmds_ch1_p, tmds_ch1_n;
    wire tmds_ch2_p, tmds_ch2_n;
    wire tmds_clk_p, tmds_clk_n;

    // DUT
    tmds_encoder #(
        .C_PIXEL_DATA_WIDTH (C_PIXEL_DATA_WIDTH)
    ) dut (
        .tmds_clk     (tmds_clk),
        .pixel_clk    (pixel_clk),
        .rst_n        (rst_n),
        .in_data_ch0  (in_data_ch0),
        .in_data_ch1  (in_data_ch1),
        .in_data_ch2  (in_data_ch2),
        .hsync_pix_clk(hsync_pix_clk),
        .vsync_pix_clk(vsync_pix_clk),
        .de_pix_clk   (de_pix_clk),
        .tmds_ch0_p   (tmds_ch0_p),
        .tmds_ch0_n   (tmds_ch0_n),
        .tmds_ch1_p   (tmds_ch1_p),
        .tmds_ch1_n   (tmds_ch1_n),
        .tmds_ch2_p   (tmds_ch2_p),
        .tmds_ch2_n   (tmds_ch2_n),
        .tmds_clk_p   (tmds_clk_p),
        .tmds_clk_n   (tmds_clk_n)
    );

    // Pixel clock ~100 MHz
    initial begin
        pixel_clk = 1'b0;
        forever #5 pixel_clk = ~pixel_clk;
    end

    // TMDS clock 10x faster (~1 GHz in sim)
    initial begin
        tmds_clk = 1'b0;
        forever #0.5 tmds_clk = ~tmds_clk;
    end

    integer i;

    initial begin
        // Init
        rst_n         = 1'b0;
        in_data_ch0   = 8'h00;
        in_data_ch1   = 8'h00;
        in_data_ch2   = 8'h00;
        hsync_pix_clk = 1'b1; // HSYNC/VSYNC usually high during active video for HDMI
        vsync_pix_clk = 1'b1;
        de_pix_clk    = 1'b0;

        // Reset phase
        @(posedge pixel_clk);
        rst_n = 1'b1;

        // Send some active video pixels (DE=1)
        de_pix_clk = 1'b1;

        // A few cycles of different colors
        for (i = 0; i < 16; i = i + 1) begin
            @(posedge pixel_clk);
            case (i)
                0:  begin in_data_ch0 <= 8'hFF; in_data_ch1 <= 8'h00; in_data_ch2 <= 8'h00; end // full blue
                1:  begin in_data_ch0 <= 8'h00; in_data_ch1 <= 8'hFF; in_data_ch2 <= 8'h00; end // full green
                2:  begin in_data_ch0 <= 8'h00; in_data_ch1 <= 8'h00; in_data_ch2 <= 8'hFF; end // full red
                default: begin
                        in_data_ch0 <= in_data_ch0 + 8'h11;
                        in_data_ch1 <= in_data_ch1 + 8'h22;
                        in_data_ch2 <= in_data_ch2 + 8'h33;
                    end
            endcase
        end

        // Simulating blanking interval 
        @(posedge pixel_clk);
        de_pix_clk    <= 1'b0;
        hsync_pix_clk <= 1'b0;
        vsync_pix_clk <= 1'b0;

        @(posedge pixel_clk);
        hsync_pix_clk <= 1'b1;
        vsync_pix_clk <= 1'b1;

        $display("Stopping tb_tmds_encoder simulation.");
        $finish;
    end

    // Used forver loop to monitor the values beacuse there are 2 clocks.
    initial begin
        $display("time\tde\tH\tV\tch0_p\tch1_p\tch2_p");
        forever begin
            @(posedge tmds_clk);
            $display("%0t\t%b\t%b\t%b\t0x%0d\t0x%0d\t0x%0d    ",$time, de_pix_clk, hsync_pix_clk, vsync_pix_clk,dut.shift_reg_ch0,dut.shift_reg_ch1,dut.shift_reg_ch2);
        end
    end

    initial
    begin
	$dumpfile("tb_tmds_encoder.vcd");
	$dumpon;
	$dumpvars();
    end
endmodule
//-------------------------------OUTPUT----------------------------------------
//Compiler version I-2014.03-2; Runtime version I-2014.03-2;  Dec  3 23:54 2025
//time	de	H	V	ch0_p	ch1_p	ch2_p
//1000	0	1	1	0x0	0x0	0x0    
//2000	0	1	1	0x0	0x0	0x0    
//3000	0	1	1	0x0	0x0	0x0    
//4000	0	1	1	0x0	0x0	0x0    
//5000	0	1	1	0x0	0x0	0x0    
//6000	1	1	1	0x0	0x0	0x0    
//7000	1	1	1	0x0	0x0	0x0    
//8000	1	1	1	0x0	0x0	0x0    
//9000	1	1	1	0x0	0x0	0x0    
//10000	1	1	1	0x0	0x0	0x0    
//11000	1	1	1	0x0	0x0	0x0    
//12000	1	1	1	0x0	0x0	0x0    
//13000	1	1	1	0x0	0x0	0x0    
//14000	1	1	1	0x0	0x0	0x0    
//15000	1	1	1	0x0	0x0	0x0    
//16000	1	1	1	0x256	0x256	0x256    
//17000	1	1	1	0x128	0x128	0x128    
//18000	1	1	1	0x64	0x64	0x64    
//19000	1	1	1	0x32	0x32	0x32    
//20000	1	1	1	0x16	0x16	0x16    
//21000	1	1	1	0x8	0x8	0x8    
//22000	1	1	1	0x4	0x4	0x4    
//23000	1	1	1	0x2	0x2	0x2    
//24000	1	1	1	0x1	0x1	0x1    
//25000	1	1	1	0x0	0x0	0x0    
//26000	1	1	1	0x1023	0x1023	0x1023    
//27000	1	1	1	0x511	0x511	0x511    
//28000	1	1	1	0x255	0x255	0x255    
//29000	1	1	1	0x127	0x127	0x127    
//30000	1	1	1	0x63	0x63	0x63    
//31000	1	1	1	0x31	0x31	0x31    
//32000	1	1	1	0x15	0x15	0x15    
//33000	1	1	1	0x7	0x7	0x7    
//34000	1	1	1	0x3	0x3	0x3    
//35000	1	1	1	0x1	0x1	0x1    
//36000	1	1	1	0x512	0x256	0x256    
//37000	1	1	1	0x256	0x128	0x128    
//38000	1	1	1	0x128	0x64	0x64    
//39000	1	1	1	0x64	0x32	0x32    
//40000	1	1	1	0x32	0x16	0x16    
//41000	1	1	1	0x16	0x8	0x8    
//42000	1	1	1	0x8	0x4	0x4    
//43000	1	1	1	0x4	0x2	0x2    
//44000	1	1	1	0x2	0x1	0x1    
//45000	1	1	1	0x1	0x0	0x0    
//46000	1	1	1	0x1023	0x255	0x1023    
//47000	1	1	1	0x511	0x127	0x511    
//48000	1	1	1	0x255	0x63	0x255    
//49000	1	1	1	0x127	0x31	0x127    
//50000	1	1	1	0x63	0x15	0x63    
//51000	1	1	1	0x31	0x7	0x31    
//52000	1	1	1	0x15	0x3	0x15    
//53000	1	1	1	0x7	0x1	0x7    
//54000	1	1	1	0x3	0x0	0x3    
//55000	1	1	1	0x1	0x0	0x1    
//56000	1	1	1	0x256	0x256	0x512    
//57000	1	1	1	0x128	0x128	0x256    
//58000	1	1	1	0x64	0x64	0x128    
//59000	1	1	1	0x32	0x32	0x64    
//60000	1	1	1	0x16	0x16	0x32    
//61000	1	1	1	0x8	0x8	0x16    
//62000	1	1	1	0x4	0x4	0x8    
//63000	1	1	1	0x2	0x2	0x4    
//64000	1	1	1	0x1	0x1	0x2    
//65000	1	1	1	0x0	0x0	0x1    
//66000	1	1	1	0x271	0x286	0x494    
//67000	1	1	1	0x135	0x143	0x247    
//68000	1	1	1	0x67	0x71	0x123    
//69000	1	1	1	0x33	0x35	0x61    
//70000	1	1	1	0x16	0x17	0x30    
//71000	1	1	1	0x8	0x8	0x15    
//72000	1	1	1	0x4	0x4	0x7    
//73000	1	1	1	0x2	0x2	0x3    
//74000	1	1	1	0x1	0x1	0x1    
//75000	1	1	1	0x0	0x0	0x0    
//76000	1	1	1	0x286	0x316	0x291    
//77000	1	1	1	0x143	0x158	0x145    
//78000	1	1	1	0x71	0x79	0x72    
//79000	1	1	1	0x35	0x39	0x36    
//80000	1	1	1	0x17	0x19	0x18    
//81000	1	1	1	0x8	0x9	0x9    
//82000	1	1	1	0x4	0x4	0x4    
//83000	1	1	1	0x2	0x2	0x2    
//84000	1	1	1	0x1	0x1	0x1    
//85000	1	1	1	0x0	0x0	0x0    
//86000	1	1	1	0x1006	0x631	0x887    
//87000	1	1	1	0x503	0x315	0x443    
//88000	1	1	1	0x251	0x157	0x221    
//89000	1	1	1	0x125	0x78	0x110    
//90000	1	1	1	0x62	0x39	0x55    
//91000	1	1	1	0x31	0x19	0x27    
//92000	1	1	1	0x15	0x9	0x13    
//93000	1	1	1	0x7	0x4	0x6    
//94000	1	1	1	0x3	0x2	0x3    
//95000	1	1	1	0x1	0x1	0x1    
//96000	1	1	1	0x316	0x376	0x19    
//97000	1	1	1	0x158	0x188	0x9    
//98000	1	1	1	0x79	0x94	0x4    
//99000	1	1	1	0x39	0x47	0x2    
//100000	1	1	1	0x19	0x23	0x1    
//101000	1	1	1	0x9	0x11	0x0    
//102000	1	1	1	0x4	0x5	0x0    
//103000	1	1	1	0x2	0x2	0x0    
//104000	1	1	1	0x1	0x1	0x0    
//105000	1	1	1	0x0	0x0	0x0    
//106000	1	1	1	0x307	0x563	0x767    
//107000	1	1	1	0x153	0x281	0x383    
//108000	1	1	1	0x76	0x140	0x191    
//109000	1	1	1	0x38	0x70	0x95    
//110000	1	1	1	0x19	0x35	0x47    
//111000	1	1	1	0x9	0x17	0x23    
//112000	1	1	1	0x4	0x8	0x11    
//113000	1	1	1	0x2	0x4	0x5    
//114000	1	1	1	0x1	0x2	0x2    
//115000	1	1	1	0x0	0x1	0x1    
//116000	1	1	1	0x136	0x238	0x784    
//117000	1	1	1	0x68	0x119	0x392    
//118000	1	1	1	0x34	0x59	0x196    
//119000	1	1	1	0x17	0x29	0x98    
//120000	1	1	1	0x8	0x14	0x49    
//121000	1	1	1	0x4	0x7	0x24    
//122000	1	1	1	0x2	0x3	0x12    
//123000	1	1	1	0x1	0x1	0x6    
//124000	1	1	1	0x0	0x0	0x3    
//125000	1	1	1	0x0	0x0	0x1    
//126000	1	1	1	0x632	0x527	0x803    
//127000	1	1	1	0x316	0x263	0x401    
//128000	1	1	1	0x158	0x131	0x200    
//129000	1	1	1	0x79	0x65	0x100    
//130000	1	1	1	0x39	0x32	0x50    
//131000	1	1	1	0x19	0x16	0x25    
//132000	1	1	1	0x9	0x8	0x12    
//133000	1	1	1	0x4	0x4	0x6    
//134000	1	1	1	0x2	0x2	0x3    
//135000	1	1	1	0x1	0x1	0x1    
//136000	1	1	1	0x376	0x496	0x728    
//137000	1	1	1	0x188	0x248	0x364    
//138000	1	1	1	0x94	0x124	0x182    
//139000	1	1	1	0x47	0x62	0x91    
//140000	1	1	1	0x23	0x31	0x45    
//141000	1	1	1	0x11	0x15	0x22    
//142000	1	1	1	0x5	0x7	0x11    
//143000	1	1	1	0x2	0x3	0x5    
//144000	1	1	1	0x1	0x1	0x2    
//145000	1	1	1	0x0	0x0	0x1    
//146000	1	1	1	0x375	0x494	0x531    
//147000	1	1	1	0x187	0x247	0x265    
//148000	1	1	1	0x93	0x123	0x132    
//149000	1	1	1	0x46	0x61	0x66    
//150000	1	1	1	0x23	0x30	0x33    
//151000	1	1	1	0x11	0x15	0x16    
//152000	1	1	1	0x5	0x7	0x8    
//153000	1	1	1	0x2	0x3	0x4    
//154000	1	1	1	0x1	0x1	0x2    
//155000	1	1	1	0x0	0x0	0x1    
//156000	1	1	1	0x563	0x460	0x1    
//157000	1	1	1	0x281	0x230	0x0    
//158000	1	1	1	0x140	0x115	0x0    
//159000	1	1	1	0x70	0x57	0x0    
//160000	1	1	1	0x35	0x28	0x0    
//161000	1	1	1	0x17	0x14	0x0    
//162000	1	1	1	0x8	0x7	0x0    
//163000	1	1	1	0x4	0x3	0x0    
//164000	1	1	1	0x2	0x1	0x0    
//165000	1	1	1	0x1	0x0	0x0    
//166000	1	1	1	0x572	0x647	0x1007    
//167000	1	1	1	0x286	0x323	0x503    
//168000	1	1	1	0x143	0x161	0x251    
//169000	1	1	1	0x71	0x80	0x125    
//170000	1	1	1	0x35	0x40	0x62    
//171000	1	1	1	0x17	0x20	0x31    
//172000	1	1	1	0x8	0x10	0x15    
//173000	1	1	1	0x4	0x5	0x7    
//174000	1	1	1	0x2	0x2	0x3    
//175000	1	1	1	0x1	0x1	0x1    
//176000	0	0	0	0x529	0x392	0x289    
//177000	0	0	0	0x264	0x196	0x144    
//178000	0	0	0	0x132	0x98	0x72    
//179000	0	0	0	0x66	0x49	0x36    
//180000	0	0	0	0x33	0x24	0x18    
//181000	0	0	0	0x16	0x12	0x9    
//182000	0	0	0	0x8	0x6	0x4    
//183000	0	0	0	0x4	0x3	0x2    
//184000	0	0	0	0x2	0x1	0x1    
//185000	0	0	0	0x1	0x0	0x0    
//Stopping tb_tmds_encoder simulation.
//
